//A 4-core system!
`define NUM_CORES 1
`define CORE_IDX_WIDTH 1
